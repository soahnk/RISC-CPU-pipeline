`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/30/2020 12:12:22 AM
// Design Name: 
// Module Name: InstructionMemory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module InstructionMemory(
    input [15:0]  pc,     
    output  [31:0] instruction
    );    
     reg [31:0] memory[1023:0];
    initial
    begin
    
//    General Purpose Registers
//    R0=0
//    R1= used for shifting
//    R2= Multiplicand
//    R3= Multiplier
//    R4= Sign of Multiplicand
//    R5= Sign of Multiplier
//    R6= Z and C comprator
//    R7= Sign comprator
//    R8= MSB of product EAX
//    R9= LSB of product  EBX
//    R10= Positive converter

//TEST numbers 
//positve and positive
//OP1>>R2 = 
//OP2>>R3 = 
//positive and negative
//OP1>>R2 = 0x1996C04F => 429310031(decimal) => 00_011001100101101_100000001001111
//OP2>>R3 = 0xF20538DC =>-1912944860(decimal) => 11_110010000001010_011100011011100
//product = -821246417147890660 => 0x8B65A743_E7298BE4
//R8/EAX = 0x8B65A743
//R9/EBX = 0xE7298BE4
//negative and negative
//OP1>>R2 = 
//OP2>>R3 = 


            ///////////load 1st number in R2
          memory[0] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[1] <= 32'b0100010_00010_00010_00000_00000_00000; // ADI: R2 <- R2 + 2 MSB's of Multiplicand
          memory[2] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[3] <= 32'b0110000_00010_00010_000000000001111; // LSL: R2 <- R2 << 15
          memory[4] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[5] <= 32'b1100010_00010_00010_011001100101101; // AIU: R2 <- R2 << (x) x=15 next MSBs of Multiplicand
          memory[6] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[7] <= 32'b0110000_00010_00010_000000000001111; // LSL: R2 <- R2 << 15
          memory[8] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[9] <= 32'b1100010_00010_00010_100000001001111; // AIU: R2 <- R2 + 15 LSBs of Multiplicand
          memory[10] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
            ///////////load 2nd number in R3
          memory[11] <= 32'b0100010_00011_00011_00000_00000_00011; //ADI: R3 <- R3 + 2 MSB's of Multiplier
          memory[12] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[13] <= 32'b0110000_00011_00011_000000000001111; // LSL: R3 <- R3 << 15
          memory[14] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[15] <= 32'b1100010_00011_00011_110010000001010; //AIU: R3 <- R3 << (x) x=15 next MSBs of Multiplier
          memory[16] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[17] <= 32'b0110000_00011_00011_000000000001111; // LSL: R3 <- R3 << 15
          memory[18] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[19] <= 32'b1100010_00011_00011_011100011011100; // AIU: R3 <- R3 + 15 LSBs of Multiplier
          memory[20] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
            ///////////check signs of both Multiplier and Multiplier
          memory[21] <= 32'b1100010_00111_00000_00000_00000_00001; // AIU: R7 <- R0 + 1
          memory[22] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[23] <= 32'b0110000_00111_00111_0000000000_11111; // LSL: R7 <- R7 << 31
          memory[24] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[25] <= 32'b0001000_00100_00111_00010_0000000000; // AND: R2 sign test to R4
          memory[26] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[27] <= 32'b0001000_00101_00111_00011_0000000000; // AND: R3 sign test to R5
          memory[28] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          /////////remove R2 sign bit
          memory[29] <= 32'b0100010_01010_00000_111111111111111; // ADI: R10 <- R0 + 1's
          memory[30] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[31] <= 32'b0000101_01010_01010_00111_0000000000; // SUB R10 <-R10,R7 
          memory[32] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[33] <= 32'b0001000_00010_01010_00010_0000000000; // AND R2 <-R10,R2
          memory[34] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          ////////////remove R3 sign bit
          memory[35] <= 32'b0001000_00011_01010_00011_0000000000; // AND R3 <-R10,R3
          memory[36] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          //////////////multiply
          memory[37] <= 32'b0110000_00110_00011_0000000000_11111; // LSL: R6 <- R3 << 31
          memory[38] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[39] <= 32'b0100000_00000_00110_000000000001101; // BZ:  if R6=0 PC <- (PC+1)+3 40030003
          /////if 0 skip add, goto shifting
          memory[40] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[41] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[42] <= 32'b0000010_01001_01001_00010_0000000000; //-- ADD	R9<-R9,R2
          memory[43] <= 32'b0000000_00000_00000_00000_0000000000; //NOP           
          //////shift         
          memory[44] <= 32'b0110000_00110_11111_0000000000_11111; // LSL: R6 <- R31 << 31
          memory[45] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          
          memory[46] <= 32'b0100000_00000_00110_000000000000100; // BZ:  if R6=0 PC <- (PC+1)+3
          //if no carry, skip add carry goto add MSBs
          memory[47] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[48] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[49] <= 32'b1100010_01000_01000_00000_00000_00001; // AIU: R8 <- R8 + 1
          memory[50] <= 32'b0000000_00000_00000_00000_0000000000; //NOP 
           
          /////add MSB's
          memory[51] <= 32'b0000010_01000_01000_00001_0000000000; //-- ADD	R8<-R8,R1 
          memory[52] <= 32'b0000000_00000_00000_00000_0000000000; //NOP 
          //shifting
          memory[53] <= 32'b0110000_00001_00001_0000000000_00001; // LSL: R1 <- R1 << 1
          memory[54] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          //test if R2 MSB 
          memory[55] <= 32'b0110001_00110_00010_0000000000_11111; // LSR: R6 <- R2 >> 31
          memory[56] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          
          memory[57] <= 32'b0100000_00000_00110_000000000000100; // BZ:  if R6=0 PC <- (PC+1)+3
          //BZ if R2 MSB ==0 skip R1=R1+1
          memory[58] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[59] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[60] <= 32'b1100010_00001_00001_00000_00000_00001; // AIU: R1 <- R1 + 1
          memory[61] <= 32'b0000000_00000_00000_00000_0000000000; //NOP 
          //////shift LSBs
          memory[62] <= 32'b0110000_00010_00010_0000000000_00001; // LSL: R2 <- R2 << 1
          memory[63] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          
          //////shift multiplier
          memory[64] <= 32'b0110001_00011_00011_0000000000_00001; // LSR: R3 <- R3 >> 1
          
          memory[65] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          /////if multiplicand=0 it's done 
          memory[66] <= 32'b0100000_00000_00011_000000000000100; // BZ: if R3=0 PC <- (PC+1)+2
          memory[67] <= 32'b0000000_00000_00000_00000_0000000000; //NOP          
          memory[68] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[69] <= 32'b1100001_00000_10101_000000000000000; // C2000000 JMR: PC <- R21
          memory[70] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          memory[71] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
          
          memory[72] <= 32'b0001100_00111_00100_00101_0000000000; // XOR R7 <- R4,R5
          memory[73] <= 32'b0000000_00000_00000_00000_0000000000; //NOP
    
          memory[74] <= 32'b0000010_01000_01000_00111_0000000000; //-- ADD	R8<-R8,R7 
          memory[75] <= 32'b0000000_00000_00000_00000_0000000000; //NOP 
          
    end                 
	assign	  instruction = memory[pc];
	   
endmodule
