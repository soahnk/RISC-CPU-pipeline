`ifndef _InstructionsParam_VH_
`define _InstructionsParam_VH_
parameter inst0  = 32'b0000000_00000_00000_00000_0000000000; // NOP
parameter inst1  = 32'b0000010_00001_00010_00011_0000000000; // ADD: R1 <- R2 + R3
parameter inst2  = 32'b0000101_00100_00001_00011_0000000000; // SUB: R4 <- R1 - R3
parameter inst3  = 32'b1100101_00001_00010_00011_0000000000; // SLT: if R2 < R3 then R1 = 1
parameter inst4  = 32'b0001000_00001_00010_00011_0000000000; // AND: R1 <- R2 AND R3
parameter inst5  = 32'b0001010_00001_00010_00011_0000000000; // OR:  R1 <- R2 OR R3
parameter inst6  = 32'b0001100_00001_00010_00011_0000000000; // XOR: R1 <- R2 XOR R3
parameter inst7  = 32'b0000001_00000_00100_00001_0000000000; // ST:  M[R4] <- R1
parameter inst8  = 32'b0100001_00100_00001_00000_0000000000; // LD:  R1 <- M[R4]
parameter inst9  = 32'b0100010_00001_00010__000000000000001; // ADI: R1 <- R2 + 1
parameter inst10 = 32'b0100101_00001_00010__000000000000001; // SBI: R1 <- R2 - 1
parameter inst11 = 32'b0101110_00001_00010__000000000000000; // NOT: R1 <- ~R2
parameter inst12 = 32'b0101000_00001_00010__000000000000001; // ANI: R1 <- R2 AND 000...1
parameter inst13 = 32'b0101010_00001_00010__000000000000000; // ORI: R1 <- R2 OR  000...0
parameter inst14 = 32'b0101100_00001_00010__000000000000000; // XRI: R1 <- R2 XOR 000...0
parameter inst15 = 32'b1100010_00001_00010__000000000000001; // AIU: R1 <- R2 + 1
parameter inst16 = 32'b1000101_00001_00010__000000000000001; // SIU: R1 <- R2 - 1
parameter inst17 = 32'b1000000_00011_00001__000000000000000; // MOV: R1 <- R3
parameter inst18 = 32'b0110000_00001_00010__000000000000001; // LSL: R1 <- R2 << 1
parameter inst19 = 32'b0110001_00001_00010__000000000000001; // LSR: R1 <- R2 >> 1
parameter inst20 = 32'b1100001_00000_00000__000000000000000; // JMR: PC <- R0
parameter inst21 = 32'b0100000_00000_00000__000000000000001; // BZ:  if R0=0 PC <- (PC+1)+1
parameter inst22 = 32'b1100000_00000_00000__000000000000001; // BNZ: if R0!=0 PC <- (PC+1)+1
parameter inst23 = 32'b1000100_00000_00000__000000000000001; // JMP: PC <- (PC+1)+1
parameter inst24 = 32'b0000111_00001_00000__000000000000000; // JML: PC <- (PC+1)+1, R1 <- PC+1
parameter instX  = 32'bX;
`endif